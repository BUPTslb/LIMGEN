module shift2_l1(
    input [1:0] a, // 输入a，2
    output [1:0] out // 输出sum
);

assign out = a * 2; // 逻辑左移

endmodule// 64位加法

