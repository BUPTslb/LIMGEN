entity test is
	port(
		i1:  in bit_vector(7 downto 0);
		i2:  in bit_vector(7 downto 0);
		out1: in bit_vector(7 downto 0);
		out2: in bit_vector(7 downto 0);
		clk:  in bit
	);	
end test;

architecture Behavioral of test is
signal in1:bit_vector(7 downto 0);
signal in1:bit_vector(7 downto 0);
signal A: bit_vector(7 downto 0);
signal B: bit_vector(7 downto 0);
signal C: bit_vector(7 downto 0);
signal D: bit_vector(7 downto 0);
signal E: bit_vector(7 downto 0);
signal F: bit_vector(7 downto 0);
signal G: bit_vector(7 downto 0);
signal H: bit_vector(7 downto 0);
signal I: bit_vector(7 downto 0);
signal J: bit_vector(7 downto 0);
signal K: bit_vector(7 downto 0);
signal L: bit_vector(7 downto 0);
signal M: bit_vector(7 downto 0);
signal N: bit_vector(7 downto 0);
signal O: bit_vector(7 downto 0);
signal P: bit_vector(7 downto 0);
signal Q: bit_vector(7 downto 0);
signal R: bit_vector(7 downto 0);
signal S: bit_vector(7 downto 0);
signal T: bit_vector(7 downto 0);

signal A1: bit_vector(7 downto 0);
signal B1: bit_vector(7 downto 0);
signal C1: bit_vector(7 downto 0);
signal D1: bit_vector(7 downto 0);
signal E1: bit_vector(7 downto 0);
signal F1: bit_vector(7 downto 0);
signal G1: bit_vector(7 downto 0);
signal H1: bit_vector(7 downto 0);
signal I1: bit_vector(7 downto 0);
signal J1: bit_vector(7 downto 0);
signal K1: bit_vector(7 downto 0);
signal L1: bit_vector(7 downto 0);
signal M1: bit_vector(7 downto 0);
signal N1: bit_vector(7 downto 0);
signal O1: bit_vector(7 downto 0);
signal P1: bit_vector(7 downto 0);
signal Q1: bit_vector(7 downto 0);
signal R1: bit_vector(7 downto 0);
signal S1: bit_vector(7 downto 0);
signal T1: bit_vector(7 downto 0);

signal A2: bit_vector(7 downto 0);
signal B2: bit_vector(7 downto 0);
signal C2: bit_vector(7 downto 0);
signal D2: bit_vector(7 downto 0);
signal E2: bit_vector(7 downto 0);
signal F2: bit_vector(7 downto 0);
signal G2: bit_vector(7 downto 0);
signal H2: bit_vector(7 downto 0);
signal I2: bit_vector(7 downto 0);
signal J2: bit_vector(7 downto 0);
signal K2: bit_vector(7 downto 0);
signal L2: bit_vector(7 downto 0);
signal M2: bit_vector(7 downto 0);
signal N2: bit_vector(7 downto 0);
signal O2: bit_vector(7 downto 0);
signal P2: bit_vector(7 downto 0);
signal Q2: bit_vector(7 downto 0);
signal R2: bit_vector(7 downto 0);
signal S2: bit_vector(7 downto 0);
signal T2: bit_vector(7 downto 0);

signal A3: bit_vector(7 downto 0);
signal B3: bit_vector(7 downto 0);
signal C3: bit_vector(7 downto 0);
signal D3: bit_vector(7 downto 0);
signal E3: bit_vector(7 downto 0);
signal F3: bit_vector(7 downto 0);
signal G3: bit_vector(7 downto 0);
signal H3: bit_vector(7 downto 0);
signal I3: bit_vector(7 downto 0);
signal J3: bit_vector(7 downto 0);
signal K3: bit_vector(7 downto 0);
signal L3: bit_vector(7 downto 0);
signal M3: bit_vector(7 downto 0);
signal N3: bit_vector(7 downto 0);
signal O3: bit_vector(7 downto 0);
signal P3: bit_vector(7 downto 0);
signal Q3: bit_vector(7 downto 0);
signal R3: bit_vector(7 downto 0);
signal S3: bit_vector(7 downto 0);
signal T3: bit_vector(7 downto 0);

begin
--当前只处理两个操作数的情况，多个呢？
process(clk)
begin
    i1 <= 101;
    i2 <= 010;
    in1 <= i1;
    in2 <= i2;
    A <= in1 * 2;
    B <= in1 or in2;
    C <= A xor B ;
    D <= not C;
    E <= C nor D;
    F <= D and E;
    G <= E or F;
    H <= F xor G;
    I <= G nor H;
    J <= H and I;
    K <= I or J;
    L <= J xor K;
    M <= K nor L;
    N <= L and M;
    O <= M or N;
    P <= N xor O;
    Q <= O nor P;
    R <= P and Q;
    S <= Q or R;
    T <= R xor S;
    A <= D xor B;
    B <= C xor A;
    C <= A xor B;
    D <= B xor C;
    E <= C xor D;
    F <= D xor E;
    G <= E xor F;
    H <= F xor G;
    I <= G xor H;
    J <= H xor I;
    K <= I xor J;
    L <= J xor K;
    M <= K xor L;
    N <= L xor M;
    O <= M xor N;
    P <= N xor O;
    Q <= O xor P;
    R <= P xor Q;
    S <= Q xor R;
    T <= R xor S;
    A <= C nor B;
    B <= D nor A;
    C <= A nor B;
    D <= B nor C;
    E <= C nor D;
    F <= D nor E;
    G <= E nor F;
    H <= F nor G;
    I <= G nor H;
    J <= H nor I;
    K <= I nor J;
    L <= J nor K;
    M <= K nor L;
    N <= L nor M;
    O <= M nor N;
    P <= N nor O;
    Q <= O nor P;
    R <= P nor Q;
    S <= Q nor R;
    T <= R nor S;
    C <= A and B;
    D <= B and C;
    A <= C and B;
    B <= D and A;
    C <= A and B;
    D <= B and C;
    E <= C and D;
    F <= D and E;
    G <= E and F;
    H <= F and G;
    I <= G and H;
    J <= H and I;
    K <= I and J;
    L <= J and K;
    M <= K and L;
    N <= L and M;
    O <= M and N;
    P <= N and O;
    Q <= O and P;
    R <= P and Q;
    S <= Q and R;
    T <= R and S;
    A <= C + B;
    B <= D + A;
    C <= A + B;
    D <= B + C;
    E <= C + D;
    F <= D + E;
    G <= E + F;
    H <= F + G;
    I <= G + H;
    J <= H + I;
    K <= I + J;
    L <= J + K;
    M <= K + L;
    N <= L + M;
    O <= M + N;
    P <= N + O;
    Q <= O + P;
    R <= P + Q;
    S <= Q + R;
    T <= R + S;
    A <= C or B;
    B <= D or A;
    C <= A or B;
    D <= B or C;
    E <= C or D;
    F <= D or E;
    G <= E or F;
    H <= F or G;
    I <= G or H;
    J <= H or I;
    K <= I or J;
    L <= J or K;
    M <= K or L;
    N <= L or M;
    O <= M or N;
    P <= N or O;
    Q <= O or P;
    R <= P or Q;
    S <= Q or R;
    T <= R or S;
    A <= not B;
    B <= not C;
    C <= not D;
    D <= not E;
    E <= not F;
    F <= not G;
    G <= not H;
    H <= not I;
    I <= not J;
    J <= not K;
    K <= not L;
    L <= not M;
    M <= not N;
    N <= not O;
    O <= not P;
    P <= not Q;
    Q <= not R;
    R <= not S;
    S <= not T;
    T <= not A;

    A1 <= in1 * 2;
    B1 <= in1 or in2;
    C1 <= A xor B ;
    D1 <= not C;
    E1 <= C nor D;
    F1 <= D and E;
    G1 <= E or F;
    H1 <= F xor G;
    I1 <= G nor H;
    J1 <= H and I;
    K1 <= I or J;
    L1 <= J xor K;
    M1 <= K nor L;
    N1 <= L and M;
    O1 <= M or N;
    P1 <= N xor O;
    Q1 <= O nor P;
    R1 <= P and Q;
    S1 <= Q or R;
    T1 <= R xor S;
    A1 <= D xor B;
    B1 <= C xor A;
    C1 <= A xor B;
    D1 <= B xor C;
    E1 <= C xor D;
    F1 <= D xor E;
    G1 <= E xor F;
    H1 <= F xor G;
    I1 <= G xor H;
    J1 <= H xor I;
    K1 <= I xor J;
    L1 <= J xor K;
    M1 <= K xor L;
    N1 <= L xor M;
    O1 <= M xor N;
    P1 <= N xor O;
    Q1 <= O xor P;
    R1 <= P xor Q;
    S1 <= Q xor R;
    T1 <= R xor S;
    A1 <= C nor B;
    B1 <= D nor A;
    C1 <= A nor B;
    D1 <= B nor C;
    E1 <= C nor D;
    F1 <= D nor E;
    G1 <= E nor F;
    H1 <= F nor G;
    I1 <= G nor H;
    J1 <= H nor I;
    K1 <= I nor J;
    L1 <= J nor K;
    M1 <= K nor L;
    N1 <= L nor M;
    O1 <= M nor N;
    P1 <= N nor O;
    Q1 <= O nor P;
    R1 <= P nor Q;
    S1 <= Q nor R;
    T1 <= R nor S;
    C1 <= A and B;
    D1 <= B and C;
    A1 <= C and B;
    B1 <= D and A;
    C1 <= A and B;
    D1 <= B and C;
    E1 <= C and D;
    F1 <= D and E;
    G1 <= E and F;
    H1 <= F and G;
    I1 <= G and H;
    J1 <= H and I;
    K1 <= I and J;
    L1 <= J and K;
    M1 <= K and L;
    N1 <= L and M;
    O1 <= M and N;
    P1 <= N and O;
    Q1 <= O and P;
    R1 <= P and Q;
    S1 <= Q and R;
    T1 <= R and S;
    A1 <= C + B;
    B1 <= D + A;
    C1 <= A + B;
    D1 <= B + C;
    E1 <= C + D;
    F1 <= D + E;
    G1 <= E + F;
    H1 <= F + G;
    I1 <= G + H;
    J1 <= H + I;
    K1 <= I + J;
    L1 <= J + K;
    M1 <= K + L;
    N1 <= L + M;
    O1 <= M + N;
    P1 <= N + O;
    Q1 <= O + P;
    R1 <= P + Q;
    S1 <= Q + R;
    T1 <= R + S;
    A1 <= C or B;
    B1 <= D or A;
    C1 <= A or B;
    D1 <= B or C;
    E1 <= C or D;
    F1 <= D or E;
    G1 <= E or F;
    H1 <= F or G;
    I1 <= G or H;
    J1 <= H or I;
    K1 <= I or J;
    L1 <= J or K;
    M1 <= K or L;
    N1 <= L or M;
    O1 <= M or N;
    P1 <= N or O;
    Q1 <= O or P;
    R1 <= P or Q;
    S1 <= Q or R;
    T1 <= R or S;
    A1 <= not B;
    B1 <= not C;
    C1 <= not D;
    D1 <= not E;
    E1 <= not F;
    F1 <= not G;
    G1 <= not H;
    H1 <= not I;
    I1 <= not J;
    J1 <= not K;
    K1 <= not L;
    L1 <= not M;
    M1 <= not N;
    N1 <= not O;
    O1 <= not P;
    P1 <= not Q;
    Q1 <= not R;
    R1 <= not S;
    S1 <= not T;
    T1 <= not A;

    A2 <= in1 * 2;
    B2 <= in1 or in2;
    C2 <= A xor B ;
    D2 <= not C;
    E2 <= C nor D;
    F2 <= D and E;
    G2 <= E or F;
    H2 <= F xor G;
    I2 <= G nor H;
    J2 <= H and I;
    K2 <= I or J;
    L2 <= J xor K;
    M2 <= K nor L;
    N2 <= L and M;
    O2 <= M or N;
    P2 <= N xor O;
    Q2 <= O nor P;
    R2 <= P and Q;
    S2 <= Q or R;
    T2 <= R xor S;
    A2 <= D xor B;
    B2 <= C xor A;
    C2 <= A xor B;
    D2 <= B xor C;
    E2 <= C xor D;
    F2 <= D xor E;
    G2 <= E xor F;
    H2 <= F xor G;
    I2 <= G xor H;
    J2 <= H xor I;
    K2 <= I xor J;
    L2 <= J xor K;
    M2 <= K xor L;
    N2 <= L xor M;
    O2 <= M xor N;
    P2 <= N xor O;
    Q2 <= O xor P;
    R2 <= P xor Q;
    S2 <= Q xor R;
    T2 <= R xor S;
    A2 <= C nor B;
    B2 <= D nor A;
    C2 <= A nor B;
    D2 <= B nor C;
    E2 <= C nor D;
    F2 <= D nor E;
    G2 <= E nor F;
    H2 <= F nor G;
    I2 <= G nor H;
    J2 <= H nor I;
    K2 <= I nor J;
    L2 <= J nor K;
    M2 <= K nor L;
    N2 <= L nor M;
    O2 <= M nor N;
    P2 <= N nor O;
    Q2 <= O nor P;
    R2 <= P nor Q;
    S2 <= Q nor R;
    T2 <= R nor S;
    C2 <= A and B;
    D2 <= B and C;
    A2 <= C and B;
    B2 <= D and A;
    C2 <= A and B;
    D2 <= B and C;
    E2 <= C and D;
    F2 <= D and E;
    G2 <= E and F;
    H2 <= F and G;
    I2 <= G and H;
    J2 <= H and I;
    K2 <= I and J;
    L2 <= J and K;
    M2 <= K and L;
    N2 <= L and M;
    O2 <= M and N;
    P2 <= N and O;
    Q2 <= O and P;
    R2 <= P and Q;
    S2 <= Q and R;
    T2 <= R and S;
    A2 <= C + B;
    B2 <= D + A;
    C2 <= A + B;
    D2 <= B + C;
    E2 <= C + D;
    F2 <= D + E;
    G2 <= E + F;
    H2 <= F + G;
    I2 <= G + H;
    J2 <= H + I;
    K2 <= I + J;
    L2 <= J + K;
    M2 <= K + L;
    N2 <= L + M;
    O2 <= M + N;
    P2 <= N + O;
    Q2 <= O + P;
    R2 <= P + Q;
    S2 <= Q + R;
    T2 <= R + S;
    A2 <= C or B;
    B2 <= D or A;
    C2 <= A or B;
    D2 <= B or C;
    E2 <= C or D;
    F2 <= D or E;
    G2 <= E or F;
    H2 <= F or G;
    I2 <= G or H;
    J2 <= H or I;
    K2 <= I or J;
    L2 <= J or K;
    M2 <= K or L;
    N2 <= L or M;
    O2 <= M or N;
    P2 <= N or O;
    Q2 <= O or P;
    R2 <= P or Q;
    S2 <= Q or R;
    T2 <= R or S;
    A2 <= not B;
    B2 <= not C;
    C2 <= not D;
    D2 <= not E;
    E2 <= not F;
    F2 <= not G;
    G2 <= not H;
    H2 <= not I;
    I2 <= not J;
    J2 <= not K;
    K2 <= not L;
    L2 <= not M;
    M2 <= not N;
    N2 <= not O;
    O2 <= not P;
    P2 <= not Q;
    Q2 <= not R;
    R2 <= not S;
    S2 <= not T;
    T2 <= not A;


    A2 <= D1 xor B1;
    B2 <= C1 xor A1;
    C2 <= A1 xor B1;
    D2 <= B1 xor C1;
    E2 <= C1 xor D1;
    F2 <= D1 xor E1;
    G2 <= E1 xor F1;
    H2 <= F1 xor G1;
    I2 <= G1 xor H1;
    J2 <= H1 xor I1;
    K2 <= I1 xor J1;
    L2 <= J1 xor K1;
    M2 <= K1 xor L1;
    N2 <= L1 xor M1;
    O2 <= M1 xor N1;
    P2 <= N1 xor O1;
    Q2 <= O1 xor P1;
    R2 <= P1 xor Q1;
    S2 <= Q1 xor R1;
    T2 <= R1 xor S1;
    A2 <= C1 nor B1;
    B2 <= D1 nor A1;
    C2 <= A1 nor B1;
    D2 <= B1 nor C1;
    E2 <= C1 nor D1;
    F2 <= D1 nor E1;
    G2 <= E1 nor F1;
    H2 <= F1 nor G1;
    I2 <= G1 nor H1;
    J2 <= H1 nor I1;
    K2 <= I1 nor J1;
    L2 <= J1 nor K1;
    M2 <= K1 nor L1;
    N2 <= L1 nor M1;
    O2 <= M1 nor N1;
    P2 <= N1 nor O1;
    Q2 <= O1 nor P1;
    R2 <= P1 nor Q1;
    S2 <= Q1 nor R1;
    T2 <= R1 nor S1;
    C2 <= A1 and B1;
    D2 <= B1 and C1;
    A2 <= C1 and B1;
    B2 <= D1 and A1;
    C2 <= A1 and B1;
    D2 <= B1 and C1;
    E2 <= C1 and D1;
    F2 <= D1 and E1;
    G2 <= E1 and F1;
    H2 <= F1 and G1;
    I2 <= G1 and H1;
    J2 <= H1 and I1;
    K2 <= I1 and J1;
    L2 <= J1 and K1;
    M2 <= K1 and L1;
    N2 <= L1 and M1;
    O2 <= M1 and N1;
    P2 <= N1 and O1;
    Q2 <= O1 and P1;
    R2 <= P1 and Q1;
    S2 <= Q1 and R1;
    T2 <= R1 and S1;
    A2 <= C1 + B1;
    B2 <= D1 + A1;
    C2 <= A1 + B1;
    D2 <= B1 + C1;
    E2 <= C1 + D1;
    F2 <= D1 + E1;
    G2 <= E1 + F1;
    H2 <= F1 + G1;
    I2 <= G1 + H1;
    J2 <= H1 + I1;
    K2 <= I1 + J1;
    L2 <= J1 + K1;
    M2 <= K1 + L1;
    N2 <= L1 + M1;
    O2 <= M1 + N1;
    P2 <= N1 + O1;
    Q2 <= O1 + P1;
    R2 <= P1 + Q1;
    S2 <= Q1 + R1;
    T2 <= R1 + S1;
    A2 <= C1 or B1;
    B2 <= D1 or A1;
    C2 <= A1 or B1;
    D2 <= B1 or C1;
    E2 <= C1 or D1;
    F2 <= D1 or E1;
    G2 <= E1 or F1;
    H2 <= F1 or G1;
    I2 <= G1 or H1;
    J2 <= H1 or I1;
    K2 <= I1 or J1;
    L2 <= J1 or K1;
    M2 <= K1 or L1;
    N2 <= L1 or M1;
    O2 <= M1 or N1;
    P2 <= N1 or O1;
    Q2 <= O1 or P1;
    R2 <= P1 or Q1;
    S2 <= Q1 or R1;
    T2 <= R1 or S1;
    A2 <= not B1;
    B2 <= not C1;
    C2 <= not D1;
    D2 <= not E1;
    E2 <= not F1;
    F2 <= not G1;
    G2 <= not H1;
    H2 <= not I1;
    I2 <= not J1;
    J2 <= not K1;
    K2 <= not L1;
    L2 <= not M1;
    M2 <= not N1;
    N2 <= not O1;
    O2 <= not P1;
    P2 <= not Q1;
    Q2 <= not R1;
    R2 <= not S1;
    S2 <= not T1;
    T2 <= not A1;

    A3 <= D2 xor B2;
    B3 <= A2 xor C2;
    C3 <= B2 xor D2;
    D3 <= C2 xor A2;
    E3 <= D2 nor B2;
    F3 <= A2 nor C2;
    G3 <= B2 nor D2;
    H3 <= C2 nor A2;
    I3 <= D2 and B2;
    J3 <= A2 and C2;
    K3 <= B2 and D2;
    L3 <= C2 and A2;
    M3 <= D2 + B2;
    N3 <= A2 + C2;
    O3 <= B2 + D2;
    P3 <= C2 + A2;
    Q3 <= D2 or B2;
    R3 <= A2 or C2;
    S3 <= B2 or D2;
    T3 <= C2 or A2;
    A3 <= D2 + B2;
    B3 <= A2 + C2;
    C3 <= B2 + D2;
    D3 <= C2 + A2;
    E3 <= D2 or B2;
    F3 <= A2 or C2;
    G3 <= B2 or D2;
    H3 <= C2 or A2;
    I3 <= D2 and B2;
    J3 <= A2 and C2;
    K3 <= B2 and D2;
    L3 <= C2 and A2;
    M3 <= D2 xor B2;
    N3 <= A2 xor C2;
    O3 <= B2 xor D2;
    P3 <= C2 xor A2;
    Q3 <= D2 nor B2;
    R3 <= A2 nor C2;
    S3 <= B2 nor D2;
    T3 <= C2 nor A2;
    A3 <= D2 and B2;
    B3 <= A2 and C2;
    C3 <= B2 and D2;
    D3 <= C2 and A2;
    E3 <= D2 xor B2;
    F3 <= A2 xor C2;
    G3 <= B2 xor D2;
    H3 <= C2 xor A2;
    I3 <= D2 nor B2;
    J3 <= A2 nor C2;
    K3 <= B2 nor D2;
    L3 <= C2 nor A2;
    M3 <= D2 or B2;
    N3 <= A2 or C2;
    O3 <= B2 or D2;
    P3 <= C2 or A2;
    Q3 <= D2 + B2;
    R3 <= A2 + C2;
    S3 <= B2 + D2;
    T3 <= C2 + A2;
    A3 <= D2 nor B2;
    B3 <= A2 nor C2;
    C3 <= B2 nor D2;
    D3 <= C2 nor A2;
    E3 <= D2 and B2;
    F3 <= A2 and C2;
    G3 <= B2 and D2;
    H3 <= C2 and A2;
    I3 <= D2 xor B2;
    J3 <= A2 xor C2;
    K3 <= B2 xor D2;
    L3 <= C2 xor A2;
    M3 <= D2 or B2;
    N3 <= A2 or C2;
    O3 <= B2 or D2;
    P3 <= C2 or A2;
    Q3 <= D2 and B2;
    R3 <= A2 and C2;
    S3 <= B2 and D2;
    T3 <= C2 and A2;





--有elseif的当前不太会处理
	if   A1<0    then
		A1 <= not A1;
	end if;

	if   B1=0    then
    	B1 <= not B1;
    end if;

	while A1<0 loop
	    A1 <= A1 xor 1;
	end loop;

--嵌套
	while D1 >0 loop
	    if D1 < 5 then
	        if A1 >0 then
	            D1<=D1+A1;
	        end if;
	    end if;

		D1 <= not D1 ;
	end loop ; -- identifier


	out1 <=A1 nor C2 ;
	out1 <=B1 nor out1;
	out1 <=C2 nor out1;
    out1 <=D1 nor out1;
    out1 <=E2 nor out1;
    out1 <=F1 nor out1;
    out1 <=G2 nor out1;
    out1 <=H1 nor out1;
    out1 <=I2 nor out1;
    out1 <=J1 nor out1;
    out1 <=K2 nor out1;
    out1 <=L1 nor out1;
    out1 <=M2 nor out1;
    out1 <=N1 nor out1;
    out1 <=O2 nor out1;
    out1 <=P1 nor out1;
    out1 <=Q2 nor out1;
    out1 <=R1 nor out1;
    out1 <=S2 nor out1;
    out1 <=T1 nor out1;

	out2 <=B1 xor D1;
	out2 <=C1 xor out2;
	out2 <=D2 xor out2;
	out2 <=E1 xor out2;
    out2 <=F2 xor out2;
    out2 <=G1 xor out2;
    out2 <=H2 xor out2;
    out2 <=I1 xor out2;
    out2 <=J2 xor out2;
    out2 <=K1 xor out2;
    out2 <=L2 xor out2;
    out2 <=M1 xor out2;
    out2 <=N2 xor out2;
    out2 <=O1 xor out2;
    out2 <=P2 xor out2;
    out2 <=Q1 xor out2;
    out2 <=R2 xor out2;
    out2 <=S1 xor out2;
    out2 <=T2 xor out2;
    out1 <=out2 xor A1;
    out2 <=out1 xor B2;
    out1 <=out2 xor C1;
    out2 <=out1 xor D2;
    out1 <=out2 xor E1;
    out2 <=out1 xor F2;
    out1 <=out2 xor G1;
    out2 <=out1 xor H2;
    out1 <=out2 xor I1;
    out2 <=out1 xor J2;
    out1 <=out2 xor K1;
    out2 <=out1 xor L2;
    out1 <=out2 xor M1;
    out2 <=out1 xor N2;
    out1 <=out2 xor O1;
    out2 <=out1 xor P2;
    out1 <=out2 xor Q1;
    out2 <=out1 xor R2;
    out1 <=out2 xor S1;
    out2 <=out1 xor T2;
    out1 <= not out2;
    out2 <= not out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;
    out1 <= out1 xor out2;
    out2 <= out2 xor out1;

end process;

end Behavioral;