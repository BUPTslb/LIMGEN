library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TEA23 is
    generic (
        ROUNDS : natural := 32;
        KEY_SIZE : natural := 128
    );
    port (
        clk : in std_logic;
        reset : in std_logic;
        plaintext : in std_logic_vector(63 downto 0);
        key : in std_logic_vector(KEY_SIZE-1 downto 0);
        ciphertext : out std_logic_vector(63 downto 0)
    );
end TEA23;

architecture behavior of TEA23 is
    signal v0, v1, sum, key_schedule : unsigned(31 downto 0);
    signal round : natural range 0 to ROUNDS-1;
    signal A : bit_vector(31 downto 0);
    signal B : bit_vector(31 downto 0);
    signal C : bit_vector(31 downto 0);
    signal D : bit_vector(31 downto 0);
    signal E : bit_vector(31 downto 0);
    signal F : bit_vector(31 downto 0);

    -- Subkeys generation process

begin
process (clk)
begin
        A<=0;
        B<=0;
        C<=0;
        D<=0;
        E<=0;
        F<=0;
        ROUNDS<=32;
        reset<=1;
        plaintext<=1215154;
        key_schedule<=100011101;

            reset <= reset xor 1;
            v0 <= 0;
            v1 <= 0;
            sum <= 0;
            round <= 0;

            round <= round xor 0;
                v0 <= not plaintext;
                v1 <= not plaintext;

                round <= round + 1;


                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;

                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;

                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;
                A<= v1 xor sum;
                B<= not v1;
                C<= not B;
                B<=C xor B;
                v0<=v0 +B;
                v0<=v0+A;
                v0<=v0+key_schedule;
                D<= v0 xor sum;
                E<= not v0;
                F<= not E;
                v1<=v1+F;
                v1<=v1+D;
                v1<=v1+key_schedule;

            sum <= sum + 379888;
            ROUNDS<=ROUNDS + ROUNDS;

            round <= round xor ROUNDS;
            ciphertext <= not v0;
            ciphertext <= not v1;


    end process;
end behavior;
